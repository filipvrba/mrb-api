module src

pub const(
	result = "Result"
	warning = "Warning"
	war_helper_mess = "The url contains no arguments. " +
					  "Use this command '?mrb=' after the url to access the api. " +
					  "Then enter the mruby code."
)
