module src

pub const(
	result = "Result"
	warning = "Warning"
	error = "Error"
	war_helper_mess = "The url contains no arguments. " +
					  "Use this command '?mrb=' after the url to access the api. " +
					  "Then enter the mruby code."
	err_token_mess_a = "Not inserted is the API Token. " +
						"Please place it after the command '?token='."
	err_token_mess_b = "Please use another token because this one is invalid."
)
